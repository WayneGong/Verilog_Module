//---------------------------------------------------------------------------
//--	文件名		:	key_in_Module.v
//--	描述		:	按键消抖模块1,按下时为低有效
//---------------------------------------------------------------------------
module key_Module
#(
	KEY_NUM	=	3
)
(
	clk,
	rst_n,
	key_in,

	key_out
);  
 
//---------------------------------------------------------------------------
//--	外部端口声明
//---------------------------------------------------------------------------
input					clk;				//时钟的端口,开发板用的50MHz晶振
input					rst_n;				//复位的端口,低电平复位
input		[ KEY_NUM-1:0]		key_in;					//对应开发板上的key_in
output		[ KEY_NUM-1:0]		key_out;				//对应开发板上的LED

//---------------------------------------------------------------------------
//--	内部端口声明
//---------------------------------------------------------------------------

reg		[31:0]			time_cnt;			//用来计数按键延迟的定时计数器
reg		[ KEY_NUM-1:0]	key_out_reg;

//设置定时器的时间为20ms
//按键按下时为低电平，没有按下时为高电平
//当按键的值不为全1时，则按键被按下，此时记录按键按下的时间，当计时的低24位为全1时，计时约为0.3秒，输出一次有效的按键值，直到按键松开


always @ (posedge clk, negedge rst_n)
begin
	if(!rst_n)							
		time_cnt	<=	20'h0;				
	else if( key_in	!= 8'hff )		//当按键的值不为全1时，则按键被按下
		time_cnt	<=	time_cnt	+	1'b1;			
	else
		time_cnt	<=	20'h0;
end


always @ (posedge clk, negedge rst_n)
begin
	if(!rst_n)								
		key_out_reg	<=	8'h00;	
	else if( time_cnt[23:0] == 24'hff_ffff ) 
		key_out_reg	<=	~key_in;			//按下的按键为低电平，取反后输出。
	else 
		key_out_reg	<=	8'h00;	
end



assign key_out = key_out_reg;	//判断按键有没有按下

endmodule


