  `timescale 1 ns / 1 ps

module AXI_Test_M #
(
	// Parameters of Axi Master Bus Interface M00_AXI
	parameter  			C_M00_AXI_START_DATA_VALUE			= 	32'hAA000000,
	parameter  			C_M00_AXI_TARGET_SLAVE_BASE_ADDR	= 	32'h40000000,
	parameter integer 	C_M00_AXI_ADDR_WIDTH				= 	32,
	parameter integer 	C_M00_AXI_DATA_WIDTH				= 	32,
	parameter integer 	C_M00_AXI_TRANSACTIONS_NUM			= 	4
)
(
	// Ports of Axi Master Bus Interface M00_AXI
	input 	wire  								m00_axi_init_axi_txn,
	output 	wire  								m00_axi_error,
	output 	wire  								m00_axi_txn_done,
	input 	wire  								m00_axi_aclk,
	input 	wire  								m00_axi_aresetn,
	output 	wire [C_M00_AXI_ADDR_WIDTH-1 : 0] 	m00_axi_awaddr,
	output 	wire [2 : 0] 						m00_axi_awprot,
	output 	wire  								m00_axi_awvalid,
	input 	wire  								m00_axi_awready,
	output 	wire [C_M00_AXI_DATA_WIDTH-1 : 0] 	m00_axi_wdata,
	output 	wire [C_M00_AXI_DATA_WIDTH/8-1 : 0] m00_axi_wstrb,
	output 	wire 								m00_axi_wvalid,
	input 	wire 								m00_axi_wready,
	input 	wire [1 : 0] 						m00_axi_bresp,
	input 	wire 								m00_axi_bvalid,
	output 	wire 								m00_axi_bready,
	output 	wire [C_M00_AXI_ADDR_WIDTH-1 : 0] 	m00_axi_araddr,
	output 	wire [2 : 0] 						m00_axi_arprot,
	output 	wire  								m00_axi_arvalid,
	input 	wire  								m00_axi_arready,
	input 	wire [C_M00_AXI_DATA_WIDTH-1 : 0] 	m00_axi_rdata,
	input 	wire [1 : 0] 						m00_axi_rresp,
	input 	wire  								m00_axi_rvalid,
	output 	wire  								m00_axi_rready
);
// Instantiation of Axi Bus Interface M00_AXI
AXI_Test_M_v1_0_M00_AXI 
#( 
	.C_M_START_DATA_VALUE		(	C_M00_AXI_START_DATA_VALUE			),
	.C_M_TARGET_SLAVE_BASE_ADDR	(	C_M00_AXI_TARGET_SLAVE_BASE_ADDR	),
	.C_M_AXI_ADDR_WIDTH			(	C_M00_AXI_ADDR_WIDTH				),
	.C_M_AXI_DATA_WIDTH			(	C_M00_AXI_DATA_WIDTH				),
	.C_M_TRANSACTIONS_NUM		(	C_M00_AXI_TRANSACTIONS_NUM			)
) AXI_Test_v1_0_M00_AXI_inst 

(
	.INIT_AXI_TXN		(	m00_axi_init_axi_txn	),
	.ERROR				(	m00_axi_error			),
	.TXN_DONE			(	m00_axi_txn_done		),
	.M_AXI_ACLK			(	m00_axi_aclk			),
	.M_AXI_ARESETN		(	m00_axi_aresetn			),
	
	.M_AXI_AW_ADDR		(	m00_axi_awaddr			),
	.M_AXI_AW_PROT		(	m00_axi_awprot			),
	.M_AXI_AW_VALID		(	m00_axi_awvalid			),
	.M_AXI_AW_READY		(	m00_axi_awready			),
	
	.M_AXI_W_DATA		(	m00_axi_wdata			),
	.M_AXI_W_STRB		(	m00_axi_wstrb			),
	.M_AXI_W_VALID		(	m00_axi_wvalid			),
	.M_AXI_W_READY		(	m00_axi_wready			),
	
	.M_AXI_B_RESP		(	m00_axi_bresp			),
	.M_AXI_B_VALID		(	m00_axi_bvalid			),
	.M_AXI_B_READY		(	m00_axi_bready			),
	
	.M_AXI_AR_ADDR		(	m00_axi_araddr			),
	.M_AXI_AR_PROT		(	m00_axi_arprot			),
	.M_AXI_AR_VALID		(	m00_axi_arvalid			),
	.M_AXI_AR_READY		(	m00_axi_arready			),
	
	.M_AXI_R_DATA		(	m00_axi_rdata			),
	.M_AXI_R_RESP		(	m00_axi_rresp			),
	.M_AXI_R_VALID		(	m00_axi_rvalid			),
	.M_AXI_R_READY		(	m00_axi_rready			)
);

// Add user logic here

// User logic ends

endmodule
